`timescale 1ns / 1ps

`include "adder.v"
`include "alu.v"
`include "controller.v"
`include "data_memory.v"
`include "inst_rom.v"
`include "mux.v"
`include "register.v"
`include "sign_extend.v"

module processor(clk, reset, serial_in, serial_valid_in, serial_ready_in, serial_rden_out, serial_out, serial_wren_out);


endmodule
