module mux #(parameter size = 1) (
  input select,
  input [size - 1:0] in_0,
  input [size - 1:0] in_1,
  output [size - 1:0] out
);

  assign out = (select) ? in_1 : in_0;

endmodule

